module processor (
  input clock,
  input rst
);

endmodule